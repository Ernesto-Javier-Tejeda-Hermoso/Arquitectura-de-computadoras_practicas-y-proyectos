//1. Definicion del modulo y sus entradas y salidas
module _and (input A, input B, output C);
//2. declarar señales/elementos internos
//NO aplica en este ejemplo
//3. Comportamiento del modulo 
//(asignaciones, instancias, conexiones)
assign C = A&B;


endmodule
